module contador ( 
	clk,
	reset,
	salida_IBV
	) ;

input  clk;
input  reset;
inout [7:0] salida_IBV;
