module comparador ( 
	a,
	b,
	c,
	d,
	eq,
	lt,
	gt
	) ;

input  a;
input  b;
input  c;
input  d;
inout  eq;
inout  lt;
inout  gt;
