module half_adder ( 
	a,
	b,
	s,
	c
	) ;

input  a;
input  b;
inout  s;
inout  c;
