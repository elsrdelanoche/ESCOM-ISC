module restador ( 
	a,
	b,
	r,
	carry
	) ;

input  a;
input  b;
inout  r;
inout  carry;
