module sumadorrestador ( 
	a,
	b,
	carry,
	estado,
	sum,
	cout
	) ;

input  a;
input  b;
input  carry;
input  estado;
inout  sum;
inout  cout;
