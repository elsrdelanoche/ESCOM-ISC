module mediosumador ( 
	a,
	b,
	sum,
	cout
	) ;

input  a;
input  b;
inout  sum;
inout  cout;
