module pines ( 
	p,
	clk,
	load,
	q
	) ;

input [3:0] p;
input  clk;
input  load;
inout [3:0] q;
