module full_adder_3bit ( 
	a,
	b,
	c_in,
	sum,
	c_out
	) ;

input [2:0] a;
input [2:0] b;
input  c_in;
inout [2:0] sum;
inout  c_out;
