module variables ( 
	a,
	y
	) ;

input  a;
inout  y;
