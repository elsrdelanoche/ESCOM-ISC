module sum_diff_2bit ( 
	a,
	b,
	operation,
	seg
	) ;

input [1:0] a;
input [1:0] b;
input  operation;
inout [6:0] seg;
