module bcd_7seg ( 
	b0,
	b1,
	b2,
	b3,
	a,
	b,
	c,
	d,
	e,
	f,
	g
	) ;

input  b0;
input  b1;
input  b2;
input  b3;
inout  a;
inout  b;
inout  c;
inout  d;
inout  e;
inout  f;
inout  g;
