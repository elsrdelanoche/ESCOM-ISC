module sumadorcompleto ( 
	a,
	b,
	carry,
	sum,
	cout
	) ;

input  a;
input  b;
input  carry;
inout  sum;
inout  cout;
