module sumador ( 
	a,
	b,
	cin,
	cout,
	s
	) ;

input  a;
input  b;
input  cin;
inout  cout;
inout  s;
